`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 15.12.2023 13:06:03
// Design Name: 
// Module Name: imageProcessingModule
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module imageProcessingModule(
input   axi_clk,
input   axi_reset_n,
//slave interface
input   i_data_valid,
input [7:0] i_data,
output  o_data_ready,
//master interface
output  o_data_valid,
output [7:0] o_data,
input   i_data_ready,
//interrupt
output  o_intr
    );
    
    wire [71:0] pixel_data;
    wire pixel_data_valid;
    wire axis_prog_full;
    wire [7:0] convolved_data;
    wire convolved_data_valid;
    
    assign o_data_ready = !axis_prog_full;
    
    imageSourceControl ISC(
        .i_clk(axi_clk),
        .i_rst(!axi_reset_n),
        .i_pixel_data(i_data),
        .i_pixel_data_valid(i_data_valid),
        .o_pixel_data(pixel_data),
        .o_pixel_data_valid(pixel_data_valid),
        .o_intr(o_intr)
    );
    
    convModule conv(
        .i_clk(axi_clk),
        .i_incoming_pixel_data(pixel_data),
        .i_pixel_data_valid(pixel_data_valid),
        .o_convolved_data(convolved_data),
        .o_convolved_data_valid(convolved_data_valid)
    );
    
    outputBuffer OB(
       .wr_rst_busy(),        // output wire wr_rst_busy
       .rd_rst_busy(),        // output wire rd_rst_busy
       .s_aclk(axi_clk),                  // input wire s_aclk
       .s_aresetn(axi_reset_n),            // input wire s_aresetn
       .s_axis_tvalid(convolved_data_valid),    // input wire s_axis_tvalid
       .s_axis_tready(),    // output wire s_axis_tready
       .s_axis_tdata(convolved_data),      // input wire [7 : 0] s_axis_tdata
       .m_axis_tvalid(o_data_valid),    // output wire m_axis_tvalid
       .m_axis_tready(i_data_ready),    // input wire m_axis_tready
       .m_axis_tdata(o_data),      // output wire [7 : 0] m_axis_tdata
       .axis_prog_full(axis_prog_full)  // output wire axis_prog_full
    );
    
endmodule
